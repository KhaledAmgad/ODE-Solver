module FixedPoint_Division_Baseline_TB#(parameter WIDTH = 16)();
  reg  [WIDTH-1:0]a,b;
  wire [WIDTH-1:0]sum;
  wire overflowFlag;
  localparam sf = 2.0**-7.0; //  scaling factor is first 7 bits 
  localparam sfUP = 2.0**7.0; //  scaling factor is first 7 bits 
  integer i,j,intSum,intA,intB;
  FixedPoint_Division_Baseline b1(a,b,sum,overflowFlag);


  initial begin
		
	
      $display("test Cases for addition Generated by loops !!");

	  for(i=0;i<65535;i=i+100) begin
            for(j=0;j<65535;j=j+100) begin
                 assign a = i;
                 assign b = j;
				 assign intA=$signed (a)*sfUP;
				 assign intB=$signed (b);
				 
				 
				 assign intSum=(intA / intB);
                 #10;
				  if($signed (sum)==$signed (intSum) && overflowFlag==0)
					$display("(Loop )%f / %f = %f, overflowFlag = %f",  $signed(a)*sf,$signed (b)*sf,$signed (sum)*sf,(overflowFlag));				
				  else
					$display("wrong (Loop ) %f / %f = %f, overflowFlag = %f,  intSum= %f ",  $signed(a)*sf,$signed (b)*sf,$signed (sum)*sf,(overflowFlag),$signed (intSum)*sf);
					

            end  
      end
	  
	  
	  
    end

  


endmodule